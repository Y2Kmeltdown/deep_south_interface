// tg_top0_1.v

// Generated using ACDS version 19.4 64

`timescale 1 ps / 1 ps
module tg_top0_1 (
		input  wire         wmc_clk_in,          //  wmc_clk_in.clk
		input  wire         wmcrst_n_in,         // wmcrst_n_in.reset_n
		input  wire         ninit_done,          //  ninit_done.ninit_done
		output wire [8:0]   awid,                //         axi.awid
		output wire [28:0]  awaddr,              //            .awaddr
		output wire [7:0]   awlen,               //            .awlen
		output wire [2:0]   awsize,              //            .awsize
		output wire [1:0]   awburst,             //            .awburst
		output wire [2:0]   awprot,              //            .awprot
		output wire [3:0]   awqos,               //            .awqos
		output wire [0:0]   awuser_ap,           //            .awuser
		output wire         awvalid,             //            .awvalid
		input  wire         awready,             //            .awready
		output wire [255:0] wdata,               //            .wdata
		output wire [31:0]  wstrb,               //            .wstrb
		output wire         wlast,               //            .wlast
		output wire         wvalid,              //            .wvalid
		input  wire         wready,              //            .wready
		input  wire [8:0]   bid,                 //            .bid
		input  wire [1:0]   bresp,               //            .bresp
		input  wire         bvalid,              //            .bvalid
		output wire         bready,              //            .bready
		output wire [8:0]   arid,                //            .arid
		output wire [28:0]  araddr,              //            .araddr
		output wire [7:0]   arlen,               //            .arlen
		output wire [2:0]   arsize,              //            .arsize
		output wire [1:0]   arburst,             //            .arburst
		output wire [2:0]   arprot,              //            .arprot
		output wire [3:0]   arqos,               //            .arqos
		output wire [0:0]   aruser_ap,           //            .aruser
		output wire         arvalid,             //            .arvalid
		input  wire         arready,             //            .arready
		input  wire [8:0]   rid,                 //            .rid
		input  wire [255:0] rdata,               //            .rdata
		input  wire [1:0]   rresp,               //            .rresp
		input  wire         rlast,               //            .rlast
		input  wire         rvalid,              //            .rvalid
		output wire         rready,              //            .rready
		input  wire         ruser_err_dbe,       //   axi_extra.ruser_err_dbe
		input  wire [31:0]  ruser_data,          //            .ruser_data
		output wire [31:0]  wuser_data,          //            .wuser_data
		output wire [3:0]   wuser_strb,          //            .wuser_strb
		output wire         traffic_gen_pass,    //   tg_status.traffic_gen_pass
		output wire         traffic_gen_fail,    //            .traffic_gen_fail
		output wire         traffic_gen_timeout  //            .traffic_gen_timeout
	);

	altera_hbm_tg_axi_top #(
		.DIAG_RUN_DEFAULT_PATTERN        (1),
		.DIAG_RUN_USER_STAGE             (0),
		.DIAG_RUN_REPEAT_STAGE           (0),
		.DIAG_RUN_STRESS_STAGE           (0),
		.DIAG_EFFICIENCY_MONITOR         (0),
		.DIAG_HBMC_TEST_PATTERN          (0),
		.DIAG_MIXED_TRAFFIC              (0),
		.DIAG_HBM_LFSR                   (0),
		.DIAG_TEST_RANDOM_AXI_READY      (0),
		.TG_USE_EFFICIENCY_PATTERN       (0),
		.SEED_OFFSET                     (1),
		.MMR_LINK                        (0),
		.MEGAFUNC_DEVICE_FAMILY          ("STRATIX 10"),
		.USE_BYTE_EN                     (0),
		.USE_HARD_CTRL                   (1),
		.USE_MMR_EN                      (1),
		.DIAG_WR_PAR                     (0),
		.DIAG_RD_PAR                     (0),
		.DIAG_SBE_CORRECT                (0),
		.DIAG_INFI_TG_ERR_TEST           (0),
		.WORD_ADDRESS_DIVISIBLE_BY       (2),
		.BURST_COUNT_DIVISIBLE_BY        (2),
		.BURST_LEN                       (2),
		.USER_DATA_EN                    (0),
		.USE_SIMPLE_TG                   (0),
		.TEST_DURATION                   ("MEDIUM"),
		.WORD_ADDR_WIDTH                 (24),
		.DIAG_TG_OOO_EN                  (0),
		.DIAG_TG_GENERATE_RW_IDS         (1),
		.USER_RFSH_ALL_EN                (0),
		.CORE_CLK_FREQ_MHZ               (250),
		.MEM_BANK_ADDR_WIDTH             (2),
		.MEM_ROW_ADDR_WIDTH              (14),
		.AVL_TO_DQ_WIDTH_RATIO           (4),
		.MEM_BANK_GROUP_WIDTH            (2),
		.MEM_STACK_ID_WIDTH              (1),
		.MEM_COL_ADDR_WIDTH              (5),
		.ROW_ADDR_LSB                    (9),
		.BANK_ADDR_LSB                   (7),
		.COL_ADDR_LSB                    (2),
		.BANK_GROUP_LSB                  (0),
		.STACK_ID_LSB                    (23),
		.BACKPRESSURE_LATENCY            (0),
		.PIPELINE_RRESP                  (0),
		.PIPELINE_BRESP                  (0),
		.CFG_TG_READ_COUNT               (5000),
		.CFG_TG_WRITE_COUNT              (2500),
		.CFG_TG_SEQUENCE                 ("TG_SEQUENCE_RANDOM"),
		.EFFICIENCY_FACTOR_NUM           (500),
		.EFFICIENCY_FACTOR_DEN           (600),
		.ENABLE_DATA_CHECK               (1),
		.ENABLE_TEST_MODE                (0),
		.DIAG_EFFICIENCY_TEST_MODE       (0),
		.C2P_CLK_RATIO                   (2),
		.PORT_AXI_AWID_WIDTH             (9),
		.PORT_AXI_AWADDR_WIDTH           (29),
		.PORT_AXI_AWLEN_WIDTH            (8),
		.PORT_AXI_AWSIZE_WIDTH           (3),
		.PORT_AXI_AWBURST_WIDTH          (2),
		.PORT_AXI_AWPROT_WIDTH           (3),
		.PORT_AXI_AWQOS_WIDTH            (4),
		.PORT_AXI_AWUSER_AP_WIDTH        (1),
		.PORT_AXI_WDATA_WIDTH            (256),
		.PORT_AXI_WSTRB_WIDTH            (32),
		.PORT_AXI_BID_WIDTH              (9),
		.PORT_AXI_BRESP_WIDTH            (2),
		.PORT_AXI_ARID_WIDTH             (9),
		.PORT_AXI_ARADDR_WIDTH           (29),
		.PORT_AXI_ARLEN_WIDTH            (8),
		.PORT_AXI_ARSIZE_WIDTH           (3),
		.PORT_AXI_ARBURST_WIDTH          (2),
		.PORT_AXI_ARPROT_WIDTH           (3),
		.PORT_AXI_ARQOS_WIDTH            (4),
		.PORT_AXI_ARUSER_AP_WIDTH        (1),
		.PORT_AXI_RID_WIDTH              (9),
		.PORT_AXI_RDATA_WIDTH            (256),
		.PORT_AXI_RRESP_WIDTH            (2),
		.PORT_AXI_EXTRA_RUSER_DATA_WIDTH (32),
		.PORT_AXI_EXTRA_WUSER_DATA_WIDTH (32),
		.PORT_AXI_EXTRA_WUSER_STRB_WIDTH (4),
		.PORT_TG_CFG_ADDRESS_WIDTH       (10),
		.PORT_TG_CFG_RDATA_WIDTH         (32),
		.PORT_TG_CFG_WDATA_WIDTH         (32),
		.PORT_EFFMON_CSR_ADDRESS_WIDTH   (10),
		.PORT_EFFMON_CSR_RDATA_WIDTH     (32),
		.PORT_EFFMON_CSR_WDATA_WIDTH     (32),
		.PORT_APB_PADDR_WIDTH            (16),
		.PORT_APB_PWDATA_WIDTH           (16),
		.PORT_APB_PSTRB_WIDTH            (2),
		.PORT_APB_PRDATA_WIDTH           (16)
	) tg0_1 (
		.wmc_clk_in               (wmc_clk_in),                           //   input,    width = 1,  wmc_clk_in.clk
		.wmcrst_n_in              (wmcrst_n_in),                          //   input,    width = 1, wmcrst_n_in.reset_n
		.ninit_done               (ninit_done),                           //   input,    width = 1,  ninit_done.ninit_done
		.awid                     (awid),                                 //  output,    width = 9,         axi.awid
		.awaddr                   (awaddr),                               //  output,   width = 29,            .awaddr
		.awlen                    (awlen),                                //  output,    width = 8,            .awlen
		.awsize                   (awsize),                               //  output,    width = 3,            .awsize
		.awburst                  (awburst),                              //  output,    width = 2,            .awburst
		.awprot                   (awprot),                               //  output,    width = 3,            .awprot
		.awqos                    (awqos),                                //  output,    width = 4,            .awqos
		.awuser_ap                (awuser_ap),                            //  output,    width = 1,            .awuser
		.awvalid                  (awvalid),                              //  output,    width = 1,            .awvalid
		.awready                  (awready),                              //   input,    width = 1,            .awready
		.wdata                    (wdata),                                //  output,  width = 256,            .wdata
		.wstrb                    (wstrb),                                //  output,   width = 32,            .wstrb
		.wlast                    (wlast),                                //  output,    width = 1,            .wlast
		.wvalid                   (wvalid),                               //  output,    width = 1,            .wvalid
		.wready                   (wready),                               //   input,    width = 1,            .wready
		.bid                      (bid),                                  //   input,    width = 9,            .bid
		.bresp                    (bresp),                                //   input,    width = 2,            .bresp
		.bvalid                   (bvalid),                               //   input,    width = 1,            .bvalid
		.bready                   (bready),                               //  output,    width = 1,            .bready
		.arid                     (arid),                                 //  output,    width = 9,            .arid
		.araddr                   (araddr),                               //  output,   width = 29,            .araddr
		.arlen                    (arlen),                                //  output,    width = 8,            .arlen
		.arsize                   (arsize),                               //  output,    width = 3,            .arsize
		.arburst                  (arburst),                              //  output,    width = 2,            .arburst
		.arprot                   (arprot),                               //  output,    width = 3,            .arprot
		.arqos                    (arqos),                                //  output,    width = 4,            .arqos
		.aruser_ap                (aruser_ap),                            //  output,    width = 1,            .aruser
		.arvalid                  (arvalid),                              //  output,    width = 1,            .arvalid
		.arready                  (arready),                              //   input,    width = 1,            .arready
		.rid                      (rid),                                  //   input,    width = 9,            .rid
		.rdata                    (rdata),                                //   input,  width = 256,            .rdata
		.rresp                    (rresp),                                //   input,    width = 2,            .rresp
		.rlast                    (rlast),                                //   input,    width = 1,            .rlast
		.rvalid                   (rvalid),                               //   input,    width = 1,            .rvalid
		.rready                   (rready),                               //  output,    width = 1,            .rready
		.ruser_err_dbe            (ruser_err_dbe),                        //   input,    width = 1,   axi_extra.ruser_err_dbe
		.ruser_data               (ruser_data),                           //   input,   width = 32,            .ruser_data
		.wuser_data               (wuser_data),                           //  output,   width = 32,            .wuser_data
		.wuser_strb               (wuser_strb),                           //  output,    width = 4,            .wuser_strb
		.traffic_gen_pass         (traffic_gen_pass),                     //  output,    width = 1,   tg_status.traffic_gen_pass
		.traffic_gen_fail         (traffic_gen_fail),                     //  output,    width = 1,            .traffic_gen_fail
		.traffic_gen_timeout      (traffic_gen_timeout),                  //  output,    width = 1,            .traffic_gen_timeout
		.tg_cfg_waitrequest       (),                                     // (terminated),                           
		.tg_cfg_read              (1'b0),                                 // (terminated),                           
		.tg_cfg_write             (1'b0),                                 // (terminated),                           
		.tg_cfg_address           (10'b0000000000),                       // (terminated),                           
		.tg_cfg_readdata          (),                                     // (terminated),                           
		.tg_cfg_writedata         (32'b00000000000000000000000000000000), // (terminated),                           
		.tg_cfg_readdatavalid     (),                                     // (terminated),                           
		.effmon_csr_waitrequest   (1'b0),                                 // (terminated),                           
		.effmon_csr_read          (),                                     // (terminated),                           
		.effmon_csr_write         (),                                     // (terminated),                           
		.effmon_csr_address       (),                                     // (terminated),                           
		.effmon_csr_readdata      (32'b00000000000000000000000000000000), // (terminated),                           
		.effmon_csr_writedata     (),                                     // (terminated),                           
		.effmon_csr_readdatavalid (1'b0),                                 // (terminated),                           
		.ur_paddr                 (),                                     // (terminated),                           
		.ur_psel                  (),                                     // (terminated),                           
		.ur_penable               (),                                     // (terminated),                           
		.ur_pwrite                (),                                     // (terminated),                           
		.ur_pwdata                (),                                     // (terminated),                           
		.ur_pstrb                 (),                                     // (terminated),                           
		.ur_prready               (1'b0),                                 // (terminated),                           
		.ur_prdata                (16'b0000000000000000)                  // (terminated),                           
	);

endmodule
